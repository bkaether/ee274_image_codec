module dct_top #(
    parameter BLOCK_SIZE = 8;
    parameter DCT_OUT_WIDTH = 52,
    parameter NUM_BLOCKS = 4800
) (
    ports
);
    
endmodule